1.00000000e+00, 6.86761958e-21
1.03514217e+00, 8.45672726e-21
1.07151931e+00, 1.04088888e-20
1.10917482e+00, 1.27134061e-20
1.14815362e+00, 1.56216009e-20
1.18850223e+00, 1.90904254e-20
1.23026877e+00, 2.31992707e-20
1.27350308e+00, 2.82457118e-20
1.31825674e+00, 3.42617162e-20
1.36458314e+00, 4.15150369e-20
1.41253754e+00, 5.00427794e-20
1.46217717e+00, 6.03691618e-20
1.51356125e+00, 7.26379251e-20
1.56675107e+00, 8.69859222e-20
1.62181010e+00, 1.04248145e-19
1.67880402e+00, 1.24456042e-19
1.73780083e+00, 1.48121145e-19
1.79887092e+00, 1.76395098e-19
1.86208714e+00, 2.09701050e-19
1.92752491e+00, 2.48303089e-19
1.99526231e+00, 2.93972862e-19
2.06538016e+00, 3.46709851e-19
2.13796209e+00, 4.08871516e-19
2.21309471e+00, 4.80754784e-19
2.29086765e+00, 5.63952253e-19
2.37137371e+00, 6.60529883e-19
2.45470892e+00, 7.74603922e-19
2.54097271e+00, 9.02412372e-19
2.63026799e+00, 1.05317133e-18
2.72270131e+00, 1.22453434e-18
2.81838293e+00, 1.42345906e-18
2.91742701e+00, 1.65212520e-18
3.01995172e+00, 1.91290626e-18
3.12607937e+00, 2.21411957e-18
3.23593657e+00, 2.55274231e-18
3.34965439e+00, 2.94243729e-18
3.46736850e+00, 3.38486017e-18
3.58921935e+00, 3.89233005e-18
3.71535229e+00, 4.46761448e-18
3.84591782e+00, 5.11431828e-18
3.98107171e+00, 5.85200415e-18
4.12097519e+00, 6.67715491e-18
4.26579519e+00, 7.61635146e-18
4.41570447e+00, 8.67235951e-18
4.57088190e+00, 9.85767504e-18
4.73151259e+00, 1.11780340e-17
4.89778819e+00, 1.26641323e-17
5.06990708e+00, 1.43241850e-17
5.24807460e+00, 1.61874468e-17
5.43250331e+00, 1.82516067e-17
5.62341325e+00, 2.05305418e-17
5.82103218e+00, 2.30735250e-17
6.02559586e+00, 2.59319770e-17
6.23734835e+00, 2.90029197e-17
6.45654229e+00, 3.24313964e-17
6.68343918e+00, 3.62191229e-17
6.91830971e+00, 4.03441217e-17
7.16143410e+00, 4.48820433e-17
7.41310241e+00, 4.98454291e-17
7.67361489e+00, 5.52389953e-17
7.94328235e+00, 6.10856368e-17
8.22242650e+00, 6.74251164e-17
8.51138038e+00, 7.43077606e-17
8.81048873e+00, 8.17320197e-17
9.12010839e+00, 8.97022166e-17
9.44060876e+00, 9.82916520e-17
9.77237221e+00, 1.07477736e-16
1.01157945e+01, 1.17283210e-16
1.04712855e+01, 1.27720434e-16
1.08392691e+01, 1.38815891e-16
1.12201845e+01, 1.50579746e-16
1.16144861e+01, 1.63012131e-16
1.20226443e+01, 1.76097610e-16
1.24451461e+01, 1.89812037e-16
1.28824955e+01, 2.04157016e-16
1.33352143e+01, 2.19230527e-16
1.38038426e+01, 2.34977075e-16
1.42889396e+01, 2.51159233e-16
1.47910839e+01, 2.68109583e-16
1.53108746e+01, 2.85557850e-16
1.58489319e+01, 3.03531490e-16
1.64058977e+01, 3.22060593e-16
1.69824365e+01, 3.41048332e-16
1.75792361e+01, 3.60323699e-16
1.81970086e+01, 3.79994748e-16
1.88364909e+01, 4.00079159e-16
1.94984460e+01, 4.20372246e-16
2.01836636e+01, 4.41005280e-16
2.08929613e+01, 4.61648828e-16
2.16271852e+01, 4.82455136e-16
2.23872114e+01, 5.03160904e-16
2.31739465e+01, 5.23989063e-16
2.39883292e+01, 5.44796616e-16
2.48313311e+01, 5.65220023e-16
2.57039578e+01, 5.85573177e-16
2.66072506e+01, 6.05867000e-16
2.75422870e+01, 6.25596005e-16
2.85101827e+01, 6.44997403e-16
2.95120923e+01, 6.63943877e-16
3.05492111e+01, 6.82524207e-16
3.16227766e+01, 7.00442731e-16
3.27340695e+01, 7.17736478e-16
3.38844156e+01, 7.34461072e-16
3.50751874e+01, 7.50458168e-16
3.63078055e+01, 7.65822098e-16
3.75837404e+01, 7.80458157e-16
3.89045145e+01, 7.94285699e-16
4.02717034e+01, 8.07233803e-16
4.16869383e+01, 8.19330282e-16
4.31519077e+01, 8.30590837e-16
4.46683592e+01, 8.41062442e-16
4.62381021e+01, 8.50592912e-16
4.78630092e+01, 8.59329940e-16
4.95450191e+01, 8.67000536e-16
5.12861384e+01, 8.73813759e-16
5.30884444e+01, 8.79941171e-16
5.49540874e+01, 8.84872640e-16
5.68852931e+01, 8.89087204e-16
5.88843655e+01, 8.92299175e-16
6.09536897e+01, 8.94826244e-16
6.30957344e+01, 8.96245860e-16
6.53130553e+01, 8.97056298e-16
6.76082975e+01, 8.97102641e-16
6.99841996e+01, 8.96185368e-16
7.24435960e+01, 8.94603786e-16
7.49894209e+01, 8.92177422e-16
7.76247117e+01, 8.89163366e-16
8.03526122e+01, 8.85263948e-16
8.31763771e+01, 8.80840341e-16
8.60993752e+01, 8.75664241e-16
8.91250938e+01, 8.70093192e-16
9.22571427e+01, 8.63602374e-16
9.54992586e+01, 8.56895830e-16
9.88553095e+01, 8.49450075e-16
1.02329299e+02, 8.41763683e-16
1.05925373e+02, 8.33516099e-16
1.09647820e+02, 8.24619075e-16
1.13501082e+02, 8.15520589e-16
1.17489755e+02, 8.06167118e-16
1.21618600e+02, 7.96435786e-16
1.25892541e+02, 7.86263422e-16
1.30316678e+02, 7.75921275e-16
1.34896288e+02, 7.65142403e-16
1.39636836e+02, 7.54393143e-16
1.44543977e+02, 7.43275282e-16
1.49623566e+02, 7.32041911e-16
1.54881662e+02, 7.20784497e-16
1.60324539e+02, 7.09169354e-16
1.65958691e+02, 6.97569551e-16
1.71790839e+02, 6.85894362e-16
1.77827941e+02, 6.74256771e-16
1.84077200e+02, 6.62452809e-16
1.90546072e+02, 6.50687540e-16
1.97242274e+02, 6.38970092e-16
2.04173794e+02, 6.27017859e-16
2.11348904e+02, 6.15371211e-16
2.18776162e+02, 6.03669742e-16
2.26464431e+02, 5.92107852e-16
2.34422882e+02, 5.80472876e-16
2.42661010e+02, 5.69091773e-16
2.51188643e+02, 5.57818506e-16
2.60015956e+02, 5.46560223e-16
2.69153480e+02, 5.35436500e-16
2.78612117e+02, 5.24419691e-16
2.88403150e+02, 5.13617140e-16
2.98538262e+02, 5.02907937e-16
3.09029543e+02, 4.92404924e-16
3.19889511e+02, 4.82126437e-16
3.31131121e+02, 4.71868170e-16
3.42767787e+02, 4.61911465e-16
3.54813389e+02, 4.52066756e-16
3.67282300e+02, 4.42444383e-16
3.80189396e+02, 4.33083294e-16
3.93550075e+02, 4.23826402e-16
4.07380278e+02, 4.14760252e-16
4.21696503e+02, 4.05945418e-16
4.36515832e+02, 3.97404998e-16
4.51855944e+02, 3.88994115e-16
4.67735141e+02, 3.80848576e-16
4.84172368e+02, 3.72891214e-16
5.01187234e+02, 3.65155080e-16
5.18800039e+02, 3.57549553e-16
5.37031796e+02, 3.50248060e-16
5.55904257e+02, 3.43151847e-16
5.75439937e+02, 3.36126472e-16
5.95662144e+02, 3.29469406e-16
6.16595002e+02, 3.23033879e-16
6.38263486e+02, 3.16708849e-16
6.60693448e+02, 3.10640370e-16
6.83911647e+02, 3.04770506e-16
7.07945784e+02, 2.99097767e-16
7.32824533e+02, 2.93642078e-16
7.58577575e+02, 2.88358949e-16
7.85235635e+02, 2.83305257e-16
8.12830516e+02, 2.78342103e-16
8.41395142e+02, 2.73577433e-16
8.70963590e+02, 2.69074251e-16
9.01571138e+02, 2.64683670e-16
9.33254301e+02, 2.60478491e-16
9.66050879e+02, 2.56460246e-16
1.00000000e+03, 2.52516837e-16
