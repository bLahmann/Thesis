1.00000000e+00, 1.00422708e-22
1.03514217e+00, 1.21670623e-22
1.07151931e+00, 1.47600657e-22
1.10917482e+00, 1.78035646e-22
1.14815362e+00, 2.14340853e-22
1.18850223e+00, 2.57621231e-22
1.23026877e+00, 3.09272109e-22
1.27350308e+00, 3.69381104e-22
1.31825674e+00, 4.39875416e-22
1.36458314e+00, 5.24880564e-22
1.41253754e+00, 6.23838979e-22
1.46217717e+00, 7.38580336e-22
1.51356125e+00, 8.73027929e-22
1.56675107e+00, 1.02912149e-21
1.62181010e+00, 1.21274153e-21
1.67880402e+00, 1.42518755e-21
1.73780083e+00, 1.67225087e-21
1.79887092e+00, 1.95474137e-21
1.86208714e+00, 2.28328544e-21
1.92752491e+00, 2.66371926e-21
1.99526231e+00, 3.09584044e-21
2.06538016e+00, 3.59672094e-21
2.13796209e+00, 4.16854303e-21
2.21309471e+00, 4.82378481e-21
2.29086765e+00, 5.55705166e-21
2.37137371e+00, 6.41523203e-21
2.45470892e+00, 7.36314746e-21
2.54097271e+00, 8.45040773e-21
2.63026799e+00, 9.69201671e-21
2.72270131e+00, 1.10832142e-20
2.81838293e+00, 1.26660846e-20
2.91742701e+00, 1.44310806e-20
3.01995172e+00, 1.64105521e-20
3.12607937e+00, 1.86510279e-20
3.23593657e+00, 2.11612449e-20
3.34965439e+00, 2.39510833e-20
3.46736850e+00, 2.70606765e-20
3.58921935e+00, 3.05689621e-20
3.71535229e+00, 3.44123070e-20
3.84591782e+00, 3.87066367e-20
3.98107171e+00, 4.34837361e-20
4.12097519e+00, 4.87783909e-20
4.26579519e+00, 5.46324147e-20
4.41570447e+00, 6.10787396e-20
4.57088190e+00, 6.81344616e-20
4.73151259e+00, 7.60700684e-20
4.89778819e+00, 8.46455774e-20
5.06990708e+00, 9.41017351e-20
5.24807460e+00, 1.04492460e-19
5.43250331e+00, 1.15812053e-19
5.62341325e+00, 1.28273055e-19
5.82103218e+00, 1.41887302e-19
6.02559586e+00, 1.56645064e-19
6.23734835e+00, 1.72651926e-19
6.45654229e+00, 1.90315284e-19
6.68343918e+00, 2.09165040e-19
6.91830971e+00, 2.29740419e-19
7.16143410e+00, 2.52149368e-19
7.41310241e+00, 2.76144352e-19
7.67361489e+00, 3.02386834e-19
7.94328235e+00, 3.30479788e-19
8.22242650e+00, 3.60900336e-19
8.51138038e+00, 3.93792319e-19
8.81048873e+00, 4.28950041e-19
9.12010839e+00, 4.66858468e-19
9.44060876e+00, 5.07365239e-19
9.77237221e+00, 5.51083057e-19
1.01157945e+01, 5.97850099e-19
1.04712855e+01, 6.48048339e-19
1.08392691e+01, 7.00897429e-19
1.12201845e+01, 7.58292136e-19
1.16144861e+01, 8.18799853e-19
1.20226443e+01, 8.83455140e-19
1.24451461e+01, 9.52857828e-19
1.28824955e+01, 1.02638540e-18
1.33352143e+01, 1.10388246e-18
1.38038426e+01, 1.18680594e-18
1.42889396e+01, 1.27492159e-18
1.47910839e+01, 1.36802324e-18
1.53108746e+01, 1.46668871e-18
1.58489319e+01, 1.57084597e-18
1.64058977e+01, 1.68119734e-18
1.69824365e+01, 1.79716599e-18
1.75792361e+01, 1.92067621e-18
1.81970086e+01, 2.05027306e-18
1.88364909e+01, 2.18658374e-18
1.94984460e+01, 2.32987432e-18
2.01836636e+01, 2.48152024e-18
2.08929613e+01, 2.64046067e-18
2.16271852e+01, 2.80823564e-18
2.23872114e+01, 2.98352634e-18
2.31739465e+01, 3.16701712e-18
2.39883292e+01, 3.36045468e-18
2.48313311e+01, 3.56187251e-18
2.57039578e+01, 3.77384409e-18
2.66072506e+01, 3.99517027e-18
2.75422870e+01, 4.22654581e-18
2.85101827e+01, 4.46691767e-18
2.95120923e+01, 4.72140381e-18
3.05492111e+01, 4.98514609e-18
3.16227766e+01, 5.25886182e-18
3.27340695e+01, 5.54729873e-18
3.38844156e+01, 5.84376200e-18
3.50751874e+01, 6.15785370e-18
3.63078055e+01, 6.47953169e-18
3.75837404e+01, 6.81606939e-18
3.89045145e+01, 7.16535165e-18
4.02717034e+01, 7.53138637e-18
4.16869383e+01, 7.90776356e-18
4.31519077e+01, 8.30075887e-18
4.46683592e+01, 8.70768694e-18
4.62381021e+01, 9.12859330e-18
4.78630092e+01, 9.56638187e-18
4.95450191e+01, 1.00184351e-17
5.12861384e+01, 1.04871845e-17
5.30884444e+01, 1.09710763e-17
5.49540874e+01, 1.14746858e-17
5.68852931e+01, 1.19955949e-17
5.88843655e+01, 1.25282743e-17
6.09536897e+01, 1.30818648e-17
6.30957344e+01, 1.36517690e-17
6.53130553e+01, 1.42420155e-17
6.76082975e+01, 1.48519506e-17
6.99841996e+01, 1.54804284e-17
7.24435960e+01, 1.61224845e-17
7.49894209e+01, 1.67879810e-17
7.76247117e+01, 1.74751172e-17
8.03526122e+01, 1.81786824e-17
8.31763771e+01, 1.89036714e-17
8.60993752e+01, 1.96525102e-17
8.91250938e+01, 2.04112199e-17
9.22571427e+01, 2.11992224e-17
9.54992586e+01, 2.20042486e-17
9.88553095e+01, 2.28363706e-17
1.02329299e+02, 2.36880529e-17
1.05925373e+02, 2.45542396e-17
1.09647820e+02, 2.54494982e-17
1.13501082e+02, 2.63573120e-17
1.17489755e+02, 2.73026134e-17
1.21618600e+02, 2.82565062e-17
1.25892541e+02, 2.92400632e-17
1.30316678e+02, 3.02449420e-17
1.34896288e+02, 3.12727709e-17
1.39636836e+02, 3.23182246e-17
1.44543977e+02, 3.33922201e-17
1.49623566e+02, 3.44829003e-17
1.54881662e+02, 3.56035925e-17
1.60324539e+02, 3.67447331e-17
1.65958691e+02, 3.79078894e-17
1.71790839e+02, 3.90993528e-17
1.77827941e+02, 4.03169433e-17
1.84077200e+02, 4.15498150e-17
1.90546072e+02, 4.28062604e-17
1.97242274e+02, 4.40991354e-17
2.04173794e+02, 4.54026430e-17
2.11348904e+02, 4.67426095e-17
2.18776162e+02, 4.80935776e-17
2.26464431e+02, 4.94755665e-17
2.34422882e+02, 5.08861873e-17
2.42661010e+02, 5.23162303e-17
2.51188643e+02, 5.37631695e-17
2.60015956e+02, 5.52545973e-17
2.69153480e+02, 5.67585413e-17
2.78612117e+02, 5.82933638e-17
2.88403150e+02, 5.98468581e-17
2.98538262e+02, 6.14301524e-17
3.09029543e+02, 6.30437458e-17
3.19889511e+02, 6.46815601e-17
3.31131121e+02, 6.63429045e-17
3.42767787e+02, 6.80194336e-17
3.54813389e+02, 6.97315902e-17
3.67282300e+02, 7.14693913e-17
3.80189396e+02, 7.32209729e-17
3.93550075e+02, 7.50106543e-17
4.07380278e+02, 7.68126304e-17
4.21696503e+02, 7.86484892e-17
4.36515832e+02, 8.05001508e-17
4.51855944e+02, 8.23853245e-17
4.67735141e+02, 8.42743936e-17
4.84172368e+02, 8.62002739e-17
5.01187234e+02, 8.81356525e-17
5.18800039e+02, 9.00935548e-17
5.37031796e+02, 9.20580090e-17
5.55904257e+02, 9.40430138e-17
5.75439937e+02, 9.60298527e-17
5.95662144e+02, 9.80521473e-17
6.16595002e+02, 1.00065496e-16
6.38263486e+02, 1.02080273e-16
6.60693448e+02, 1.04101096e-16
6.83911647e+02, 1.06103107e-16
7.07945784e+02, 1.08102575e-16
7.32824533e+02, 1.10088654e-16
7.58577575e+02, 1.12056377e-16
7.85235635e+02, 1.13984295e-16
8.12830516e+02, 1.15891038e-16
8.41395142e+02, 1.17780552e-16
8.70963590e+02, 1.19588490e-16
9.01571138e+02, 1.21344041e-16
9.33254301e+02, 1.23056388e-16
9.66050879e+02, 1.24695579e-16
1.00000000e+03, 1.26260902e-16
