1.00000000e+00, 2.76689318e-28
1.03514217e+00, 3.88072946e-28
1.07151931e+00, 5.45864972e-28
1.10917482e+00, 7.76365770e-28
1.14815362e+00, 1.12516688e-27
1.18850223e+00, 1.58720671e-27
1.23026877e+00, 2.24898108e-27
1.27350308e+00, 3.12263878e-27
1.31825674e+00, 4.44311180e-27
1.36458314e+00, 6.30101647e-27
1.41253754e+00, 8.79415525e-27
1.46217717e+00, 1.21595863e-26
1.51356125e+00, 1.69533780e-26
1.56675107e+00, 2.26097523e-26
1.62181010e+00, 3.13011082e-26
1.67880402e+00, 4.25391438e-26
1.73780083e+00, 5.82536632e-26
1.79887092e+00, 8.01364988e-26
1.86208714e+00, 1.07139083e-25
1.92752491e+00, 1.42954000e-25
1.99526231e+00, 1.91322808e-25
2.06538016e+00, 2.52145580e-25
2.13796209e+00, 3.35656274e-25
2.21309471e+00, 4.49043374e-25
2.29086765e+00, 5.89579408e-25
2.37137371e+00, 7.71220374e-25
2.45470892e+00, 1.00728209e-24
2.54097271e+00, 1.32258736e-24
2.63026799e+00, 1.73091557e-24
2.72270131e+00, 2.24122676e-24
2.81838293e+00, 2.90333598e-24
2.91742701e+00, 3.75625617e-24
3.01995172e+00, 4.83485375e-24
3.12607937e+00, 6.17520381e-24
3.23593657e+00, 7.89025221e-24
3.34965439e+00, 1.00066159e-23
3.46736850e+00, 1.27547190e-23
3.58921935e+00, 1.61477789e-23
3.71535229e+00, 2.02783340e-23
3.84591782e+00, 2.56848568e-23
3.98107171e+00, 3.21396040e-23
4.12097519e+00, 4.03114108e-23
4.26579519e+00, 5.02360934e-23
4.41570447e+00, 6.26896743e-23
4.57088190e+00, 7.74639301e-23
4.73151259e+00, 9.58058426e-23
4.89778819e+00, 1.18356335e-22
5.06990708e+00, 1.45735488e-22
5.24807460e+00, 1.78703485e-22
5.43250331e+00, 2.18329408e-22
5.62341325e+00, 2.67306632e-22
5.82103218e+00, 3.25950462e-22
6.02559586e+00, 3.94734612e-22
6.23734835e+00, 4.79291025e-22
6.45654229e+00, 5.80527908e-22
6.68343918e+00, 7.00811090e-22
6.91830971e+00, 8.42630659e-22
7.16143410e+00, 1.00931867e-21
7.41310241e+00, 1.20802806e-21
7.67361489e+00, 1.44394921e-21
7.94328235e+00, 1.72275905e-21
8.22242650e+00, 2.05026235e-21
8.51138038e+00, 2.43263744e-21
8.81048873e+00, 2.87371559e-21
9.12010839e+00, 3.40252743e-21
9.44060876e+00, 4.00645223e-21
9.77237221e+00, 4.71611655e-21
1.01157945e+01, 5.52849549e-21
1.04712855e+01, 6.48409304e-21
1.08392691e+01, 7.56621593e-21
1.12201845e+01, 8.82811545e-21
1.16144861e+01, 1.02886107e-20
1.20226443e+01, 1.19531133e-20
1.24451461e+01, 1.38407058e-20
1.28824955e+01, 1.60282250e-20
1.33352143e+01, 1.85013633e-20
1.38038426e+01, 2.13164506e-20
1.42889396e+01, 2.45072803e-20
1.47910839e+01, 2.81239358e-20
1.53108746e+01, 3.22866934e-20
1.58489319e+01, 3.69441092e-20
1.64058977e+01, 4.22056811e-20
1.69824365e+01, 4.80846594e-20
1.75792361e+01, 5.47186085e-20
1.81970086e+01, 6.21167508e-20
1.88364909e+01, 7.04338678e-20
1.94984460e+01, 7.98037837e-20
2.01836636e+01, 9.02162664e-20
2.08929613e+01, 1.01718879e-19
2.16271852e+01, 1.14585431e-19
2.23872114e+01, 1.28822572e-19
2.31739465e+01, 1.44727878e-19
2.39883292e+01, 1.62140248e-19
2.48313311e+01, 1.81577431e-19
2.57039578e+01, 2.02805091e-19
2.66072506e+01, 2.26415881e-19
2.75422870e+01, 2.52294795e-19
2.85101827e+01, 2.80384998e-19
2.95120923e+01, 3.11620827e-19
3.05492111e+01, 3.45700353e-19
3.16227766e+01, 3.82753157e-19
3.27340695e+01, 4.23583121e-19
3.38844156e+01, 4.67692709e-19
3.50751874e+01, 5.15830419e-19
3.63078055e+01, 5.68242524e-19
3.75837404e+01, 6.25180744e-19
3.89045145e+01, 6.86439681e-19
4.02717034e+01, 7.53543527e-19
4.16869383e+01, 8.25115653e-19
4.31519077e+01, 9.03555989e-19
4.46683592e+01, 9.87625632e-19
4.62381021e+01, 1.07767218e-18
4.78630092e+01, 1.17529278e-18
4.95450191e+01, 1.27933638e-18
5.12861384e+01, 1.39159058e-18
5.30884444e+01, 1.51144716e-18
5.49540874e+01, 1.64054635e-18
5.68852931e+01, 1.77797247e-18
5.88843655e+01, 1.92417334e-18
6.09536897e+01, 2.08013271e-18
6.30957344e+01, 2.24775099e-18
6.53130553e+01, 2.42345828e-18
6.76082975e+01, 2.61310968e-18
6.99841996e+01, 2.81343105e-18
7.24435960e+01, 3.02411091e-18
7.49894209e+01, 3.24962533e-18
7.76247117e+01, 3.48727744e-18
8.03526122e+01, 3.73894315e-18
8.31763771e+01, 4.00304707e-18
8.60993752e+01, 4.28170452e-18
8.91250938e+01, 4.57569569e-18
9.22571427e+01, 4.88502169e-18
9.54992586e+01, 5.20990311e-18
9.88553095e+01, 5.55274531e-18
1.02329299e+02, 5.90850508e-18
1.05925373e+02, 6.28378165e-18
1.09647820e+02, 6.67683588e-18
1.13501082e+02, 7.08596989e-18
1.17489755e+02, 7.51508976e-18
1.21618600e+02, 7.95948890e-18
1.25892541e+02, 8.42351941e-18
1.30316678e+02, 8.90681490e-18
1.34896288e+02, 9.40905740e-18
1.39636836e+02, 9.93152037e-18
1.44543977e+02, 1.04734596e-17
1.49623566e+02, 1.10344701e-17
1.54881662e+02, 1.16120946e-17
1.60324539e+02, 1.22113697e-17
1.65958691e+02, 1.28298898e-17
1.71790839e+02, 1.34714629e-17
1.77827941e+02, 1.41268190e-17
1.84077200e+02, 1.48041867e-17
1.90546072e+02, 1.55023294e-17
1.97242274e+02, 1.62186750e-17
2.04173794e+02, 1.69575846e-17
2.11348904e+02, 1.77084534e-17
2.18776162e+02, 1.84812474e-17
2.26464431e+02, 1.92709708e-17
2.34422882e+02, 2.00787456e-17
2.42661010e+02, 2.09044300e-17
2.51188643e+02, 2.17485350e-17
2.60015956e+02, 2.26080414e-17
2.69153480e+02, 2.34830551e-17
2.78612117e+02, 2.43803241e-17
2.88403150e+02, 2.52869971e-17
2.98538262e+02, 2.62087145e-17
3.09029543e+02, 2.71492662e-17
3.19889511e+02, 2.81022952e-17
3.31131121e+02, 2.90661392e-17
3.42767787e+02, 3.00469920e-17
3.54813389e+02, 3.10398403e-17
3.67282300e+02, 3.20465887e-17
3.80189396e+02, 3.30632250e-17
3.93550075e+02, 3.40906055e-17
4.07380278e+02, 3.51358692e-17
4.21696503e+02, 3.61848573e-17
4.36515832e+02, 3.72415971e-17
4.51855944e+02, 3.83066223e-17
4.67735141e+02, 3.93919010e-17
4.84172368e+02, 4.04772572e-17
5.01187234e+02, 4.15740068e-17
5.18800039e+02, 4.26793360e-17
5.37031796e+02, 4.37870626e-17
5.55904257e+02, 4.49001550e-17
5.75439937e+02, 4.60255119e-17
5.95662144e+02, 4.71532503e-17
6.16595002e+02, 4.82853681e-17
6.38263486e+02, 4.94248421e-17
6.60693448e+02, 5.05748746e-17
6.83911647e+02, 5.17134885e-17
7.07945784e+02, 5.28622347e-17
7.32824533e+02, 5.40205854e-17
7.58577575e+02, 5.51839437e-17
7.85235635e+02, 5.63370676e-17
8.12830516e+02, 5.74973587e-17
8.41395142e+02, 5.86568990e-17
8.70963590e+02, 5.98172804e-17
9.01571138e+02, 6.09843751e-17
9.33254301e+02, 6.21474541e-17
9.66050879e+02, 6.33107528e-17
1.00000000e+03, 6.44732849e-17
