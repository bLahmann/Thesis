1.00000000e+00, 0.00000000e+00
1.03514217e+00, 0.00000000e+00
1.07151931e+00, 0.00000000e+00
1.10917482e+00, 0.00000000e+00
1.14815362e+00, 0.00000000e+00
1.18850223e+00, 0.00000000e+00
1.23026877e+00, 1.11425029e-32
1.27350308e+00, 0.00000000e+00
1.31825674e+00, 9.05668457e-33
1.36458314e+00, 1.20957720e-32
1.41253754e+00, 4.14055969e-32
1.46217717e+00, 8.75672306e-32
1.51356125e+00, 9.07184526e-32
1.56675107e+00, 1.58532331e-31
1.62181010e+00, 4.32019182e-31
1.67880402e+00, 6.62917557e-31
1.73780083e+00, 9.15166590e-31
1.79887092e+00, 1.79724529e-30
1.86208714e+00, 2.50583785e-30
1.92752491e+00, 4.51197775e-30
1.99526231e+00, 7.83665196e-30
2.06538016e+00, 1.15099626e-29
2.13796209e+00, 1.83264860e-29
2.21309471e+00, 2.70887403e-29
2.29086765e+00, 4.56176841e-29
2.37137371e+00, 6.45256739e-29
2.45470892e+00, 9.53982260e-29
2.54097271e+00, 1.39295371e-28
2.63026799e+00, 1.97910792e-28
2.72270131e+00, 2.80368235e-28
2.81838293e+00, 4.03172469e-28
2.91742701e+00, 5.53714931e-28
3.01995172e+00, 7.61233624e-28
3.12607937e+00, 1.04485071e-27
3.23593657e+00, 1.43125674e-27
3.34965439e+00, 1.94831962e-27
3.46736850e+00, 2.57839897e-27
3.58921935e+00, 3.41798780e-27
3.71535229e+00, 4.54283971e-27
3.84591782e+00, 5.96349428e-27
3.98107171e+00, 7.82338313e-27
4.12097519e+00, 1.01350706e-26
4.26579519e+00, 1.33349020e-26
4.41570447e+00, 1.72093432e-26
4.57088190e+00, 2.21664650e-26
4.73151259e+00, 2.87370970e-26
4.89778819e+00, 3.71765840e-26
5.06990708e+00, 4.76295864e-26
5.24807460e+00, 6.19379751e-26
5.43250331e+00, 7.85463188e-26
5.62341325e+00, 1.01837917e-25
5.82103218e+00, 1.31958372e-25
6.02559586e+00, 1.68795372e-25
6.23734835e+00, 2.14944930e-25
6.45654229e+00, 2.77222387e-25
6.68343918e+00, 3.59753506e-25
6.91830971e+00, 4.65942810e-25
7.16143410e+00, 5.97940749e-25
7.41310241e+00, 7.65346090e-25
7.67361489e+00, 9.78994650e-25
7.94328235e+00, 1.25346358e-24
8.22242650e+00, 1.60915661e-24
8.51138038e+00, 2.05713245e-24
8.81048873e+00, 2.63370523e-24
9.12010839e+00, 3.36307919e-24
9.44060876e+00, 4.30579146e-24
9.77237221e+00, 5.48157673e-24
1.01157945e+01, 6.97267338e-24
1.04712855e+01, 8.82464000e-24
1.08392691e+01, 1.12415783e-23
1.12201845e+01, 1.42159517e-23
1.16144861e+01, 1.78262206e-23
1.20226443e+01, 2.24418588e-23
1.24451461e+01, 2.84495203e-23
1.28824955e+01, 3.58923545e-23
1.33352143e+01, 4.46246128e-23
1.38038426e+01, 5.60503922e-23
1.42889396e+01, 7.00122326e-23
1.47910839e+01, 8.71391048e-23
1.53108746e+01, 1.07732916e-22
1.58489319e+01, 1.33958369e-22
1.64058977e+01, 1.65973718e-22
1.69824365e+01, 2.04901851e-22
1.75792361e+01, 2.52296334e-22
1.81970086e+01, 3.10597417e-22
1.88364909e+01, 3.79632581e-22
1.94984460e+01, 4.66175561e-22
2.01836636e+01, 5.67918207e-22
2.08929613e+01, 6.93317519e-22
2.16271852e+01, 8.40178832e-22
2.23872114e+01, 1.02325496e-21
2.31739465e+01, 1.23674998e-21
2.39883292e+01, 1.49317546e-21
2.48313311e+01, 1.80062708e-21
2.57039578e+01, 2.16317604e-21
2.66072506e+01, 2.59572482e-21
2.75422870e+01, 3.10974980e-21
2.85101827e+01, 3.70733282e-21
2.95120923e+01, 4.41940440e-21
3.05492111e+01, 5.26691936e-21
3.16227766e+01, 6.24700965e-21
3.27340695e+01, 7.39540792e-21
3.38844156e+01, 8.74513451e-21
3.50751874e+01, 1.03325194e-20
3.63078055e+01, 1.21388707e-20
3.75837404e+01, 1.42594955e-20
3.89045145e+01, 1.67123716e-20
4.02717034e+01, 1.95646098e-20
4.16869383e+01, 2.28077123e-20
4.31519077e+01, 2.65863024e-20
4.46683592e+01, 3.09407344e-20
4.62381021e+01, 3.58827520e-20
4.78630092e+01, 4.14889097e-20
4.95450191e+01, 4.80552509e-20
5.12861384e+01, 5.54050640e-20
5.30884444e+01, 6.38207809e-20
5.49540874e+01, 7.33603466e-20
5.68852931e+01, 8.40625301e-20
5.88843655e+01, 9.63139010e-20
6.09536897e+01, 1.10060677e-19
6.30957344e+01, 1.25509605e-19
6.53130553e+01, 1.42733707e-19
6.76082975e+01, 1.62334513e-19
6.99841996e+01, 1.84172259e-19
7.24435960e+01, 2.08655526e-19
7.49894209e+01, 2.35766260e-19
7.76247117e+01, 2.66422903e-19
8.03526122e+01, 2.99890729e-19
8.31763771e+01, 3.37763604e-19
8.60993752e+01, 3.79210113e-19
8.91250938e+01, 4.24778321e-19
9.22571427e+01, 4.75369231e-19
9.54992586e+01, 5.31247125e-19
9.88553095e+01, 5.92567138e-19
1.02329299e+02, 6.60459571e-19
1.05925373e+02, 7.34493872e-19
1.09647820e+02, 8.15445529e-19
1.13501082e+02, 9.04087845e-19
1.17489755e+02, 1.00147335e-18
1.21618600e+02, 1.10754663e-18
1.25892541e+02, 1.22236418e-18
1.30316678e+02, 1.34688741e-18
1.34896288e+02, 1.48279936e-18
1.39636836e+02, 1.62957274e-18
1.44543977e+02, 1.78893118e-18
1.49623566e+02, 1.96191865e-18
1.54881662e+02, 2.14711083e-18
1.60324539e+02, 2.34702598e-18
1.65958691e+02, 2.56331191e-18
1.71790839e+02, 2.79544645e-18
1.77827941e+02, 3.04437801e-18
1.84077200e+02, 3.31184508e-18
1.90546072e+02, 3.59828806e-18
1.97242274e+02, 3.90537821e-18
2.04173794e+02, 4.23350204e-18
2.11348904e+02, 4.58558588e-18
2.18776162e+02, 4.95808481e-18
2.26464431e+02, 5.36066489e-18
2.34422882e+02, 5.78757623e-18
2.42661010e+02, 6.24036269e-18
2.51188643e+02, 6.72599510e-18
2.60015956e+02, 7.23873968e-18
2.69153480e+02, 7.78658195e-18
2.78612117e+02, 8.37181582e-18
2.88403150e+02, 8.98785407e-18
2.98538262e+02, 9.63731266e-18
3.09029543e+02, 1.03344525e-17
3.19889511e+02, 1.10774706e-17
3.31131121e+02, 1.18583421e-17
3.42767787e+02, 1.26892201e-17
3.54813389e+02, 1.35606039e-17
3.67282300e+02, 1.44900785e-17
3.80189396e+02, 1.54772746e-17
3.93550075e+02, 1.65119360e-17
4.07380278e+02, 1.76105598e-17
4.21696503e+02, 1.87716090e-17
4.36515832e+02, 1.99960900e-17
4.51855944e+02, 2.12876665e-17
4.67735141e+02, 2.26517174e-17
4.84172368e+02, 2.40843353e-17
5.01187234e+02, 2.55937082e-17
5.18800039e+02, 2.71813695e-17
5.37031796e+02, 2.88566917e-17
5.55904257e+02, 3.06091381e-17
5.75439937e+02, 3.24472697e-17
5.95662144e+02, 3.43723937e-17
6.16595002e+02, 3.64076055e-17
6.38263486e+02, 3.85258660e-17
6.60693448e+02, 4.07133189e-17
6.83911647e+02, 4.30227306e-17
7.07945784e+02, 4.54270203e-17
7.32824533e+02, 4.79277210e-17
7.58577575e+02, 5.05416522e-17
7.85235635e+02, 5.32527546e-17
8.12830516e+02, 5.60404506e-17
8.41395142e+02, 5.89356110e-17
8.70963590e+02, 6.19540224e-17
9.01571138e+02, 6.50606091e-17
9.33254301e+02, 6.82590277e-17
9.66050879e+02, 7.15632851e-17
1.00000000e+03, 7.49579940e-17
