1.00000000e+00, 6.61915316e-24
1.03514217e+00, 8.44359893e-24
1.07151931e+00, 1.07193463e-23
1.10917482e+00, 1.34922329e-23
1.14815362e+00, 1.69261862e-23
1.18850223e+00, 2.13479964e-23
1.23026877e+00, 2.65892936e-23
1.27350308e+00, 3.32065375e-23
1.31825674e+00, 4.13040142e-23
1.36458314e+00, 5.12474316e-23
1.41253754e+00, 6.33907769e-23
1.46217717e+00, 7.83184330e-23
1.51356125e+00, 9.61493784e-23
1.56675107e+00, 1.18249489e-22
1.62181010e+00, 1.44714626e-22
1.67880402e+00, 1.76722792e-22
1.73780083e+00, 2.15018647e-22
1.79887092e+00, 2.62020208e-22
1.86208714e+00, 3.16389254e-22
1.92752491e+00, 3.82673340e-22
1.99526231e+00, 4.62136225e-22
2.06538016e+00, 5.54405804e-22
2.13796209e+00, 6.66414259e-22
2.21309471e+00, 7.96838981e-22
2.29086765e+00, 9.51977273e-22
2.37137371e+00, 1.13154085e-21
2.45470892e+00, 1.34467983e-21
2.54097271e+00, 1.59587789e-21
2.63026799e+00, 1.88983644e-21
2.72270131e+00, 2.22971125e-21
2.81838293e+00, 2.62683898e-21
2.91742701e+00, 3.08868138e-21
3.01995172e+00, 3.61880897e-21
3.12607937e+00, 4.23955305e-21
3.23593657e+00, 4.94662495e-21
3.34965439e+00, 5.76637886e-21
3.46736850e+00, 6.71275018e-21
3.58921935e+00, 7.78410171e-21
3.71535229e+00, 9.02557039e-21
3.84591782e+00, 1.04306398e-20
3.98107171e+00, 1.20335162e-20
4.12097519e+00, 1.38602877e-20
4.26579519e+00, 1.59231874e-20
4.41570447e+00, 1.82612087e-20
4.57088190e+00, 2.09345384e-20
4.73151259e+00, 2.39369752e-20
4.89778819e+00, 2.72907075e-20
5.06990708e+00, 3.10918295e-20
5.24807460e+00, 3.53406048e-20
5.43250331e+00, 4.01402090e-20
5.62341325e+00, 4.54659448e-20
5.82103218e+00, 5.14496691e-20
6.02559586e+00, 5.81009087e-20
6.23734835e+00, 6.55114151e-20
6.45654229e+00, 7.37272430e-20
6.68343918e+00, 8.28128031e-20
6.91830971e+00, 9.29480188e-20
7.16143410e+00, 1.04155753e-19
7.41310241e+00, 1.16563173e-19
7.67361489e+00, 1.30064341e-19
7.94328235e+00, 1.45112477e-19
8.22242650e+00, 1.61548027e-19
8.51138038e+00, 1.79513646e-19
8.81048873e+00, 1.99459495e-19
9.12010839e+00, 2.21064376e-19
9.44060876e+00, 2.44686035e-19
9.77237221e+00, 2.70417069e-19
1.01157945e+01, 2.98307137e-19
1.04712855e+01, 3.28931884e-19
1.08392691e+01, 3.62007652e-19
1.12201845e+01, 3.97789284e-19
1.16144861e+01, 4.36593552e-19
1.20226443e+01, 4.78537483e-19
1.24451461e+01, 5.24010610e-19
1.28824955e+01, 5.72693373e-19
1.33352143e+01, 6.25437057e-19
1.38038426e+01, 6.81994182e-19
1.42889396e+01, 7.42173553e-19
1.47910839e+01, 8.07663373e-19
1.53108746e+01, 8.77274319e-19
1.58489319e+01, 9.51763803e-19
1.64058977e+01, 1.03082083e-18
1.69824365e+01, 1.11613403e-18
1.75792361e+01, 1.20674880e-18
1.81970086e+01, 1.30308141e-18
1.88364909e+01, 1.40489796e-18
1.94984460e+01, 1.51361203e-18
2.01836636e+01, 1.62905886e-18
2.08929613e+01, 1.75070078e-18
2.16271852e+01, 1.88001368e-18
2.23872114e+01, 2.01669274e-18
2.31739465e+01, 2.16133157e-18
2.39883292e+01, 2.31279089e-18
2.48313311e+01, 2.47322133e-18
2.57039578e+01, 2.64232444e-18
2.66072506e+01, 2.81913256e-18
2.75422870e+01, 3.00541539e-18
2.85101827e+01, 3.20157368e-18
2.95120923e+01, 3.40656962e-18
3.05492111e+01, 3.62248328e-18
3.16227766e+01, 3.84654234e-18
3.27340695e+01, 4.08173678e-18
3.38844156e+01, 4.32838305e-18
3.50751874e+01, 4.58487568e-18
3.63078055e+01, 4.85422909e-18
3.75837404e+01, 5.13345318e-18
3.89045145e+01, 5.42263225e-18
4.02717034e+01, 5.72739678e-18
4.16869383e+01, 6.04296058e-18
4.31519077e+01, 6.37145720e-18
4.46683592e+01, 6.71246575e-18
4.62381021e+01, 7.06760995e-18
4.78630092e+01, 7.43526362e-18
4.95450191e+01, 7.81694108e-18
5.12861384e+01, 8.21413864e-18
5.30884444e+01, 8.62375404e-18
5.49540874e+01, 9.04943479e-18
5.68852931e+01, 9.48791519e-18
5.88843655e+01, 9.94673653e-18
6.09536897e+01, 1.04175579e-17
6.30957344e+01, 1.09075653e-17
6.53130553e+01, 1.14128297e-17
6.76082975e+01, 1.19357287e-17
6.99841996e+01, 1.24754617e-17
7.24435960e+01, 1.30365376e-17
7.49894209e+01, 1.36126930e-17
7.76247117e+01, 1.42094661e-17
8.03526122e+01, 1.48271181e-17
8.31763771e+01, 1.54657281e-17
8.60993752e+01, 1.61293255e-17
8.91250938e+01, 1.68113821e-17
9.22571427e+01, 1.75184557e-17
9.54992586e+01, 1.82514973e-17
9.88553095e+01, 1.90068837e-17
1.02329299e+02, 1.97871093e-17
1.05925373e+02, 2.05981901e-17
1.09647820e+02, 2.14346106e-17
1.13501082e+02, 2.23027828e-17
1.17489755e+02, 2.32055332e-17
1.21618600e+02, 2.41323144e-17
1.25892541e+02, 2.50956534e-17
1.30316678e+02, 2.60970799e-17
1.34896288e+02, 2.71376319e-17
1.39636836e+02, 2.81998640e-17
1.44543977e+02, 2.93171736e-17
1.49623566e+02, 3.04687881e-17
1.54881662e+02, 3.16656844e-17
1.60324539e+02, 3.29032522e-17
1.65958691e+02, 3.41916932e-17
1.71790839e+02, 3.55147452e-17
1.77827941e+02, 3.69009908e-17
1.84077200e+02, 3.83225077e-17
1.90546072e+02, 3.98020095e-17
1.97242274e+02, 4.13188104e-17
2.04173794e+02, 4.28926219e-17
2.11348904e+02, 4.45241140e-17
2.18776162e+02, 4.62015401e-17
2.26464431e+02, 4.79256240e-17
2.34422882e+02, 4.96853822e-17
2.42661010e+02, 5.15113668e-17
2.51188643e+02, 5.33704361e-17
2.60015956e+02, 5.52895181e-17
2.69153480e+02, 5.72334994e-17
2.78612117e+02, 5.91956289e-17
2.88403150e+02, 6.12383779e-17
2.98538262e+02, 6.32897310e-17
3.09029543e+02, 6.53664249e-17
3.19889511e+02, 6.74744128e-17
3.31131121e+02, 6.95840907e-17
3.42767787e+02, 7.17164103e-17
3.54813389e+02, 7.38595664e-17
3.67282300e+02, 7.60001837e-17
3.80189396e+02, 7.81306564e-17
3.93550075e+02, 8.02675131e-17
4.07380278e+02, 8.23701293e-17
4.21696503e+02, 8.44503003e-17
4.36515832e+02, 8.65232385e-17
4.51855944e+02, 8.85336337e-17
4.67735141e+02, 9.05206756e-17
4.84172368e+02, 9.24441132e-17
5.01187234e+02, 9.43266911e-17
5.18800039e+02, 9.61454445e-17
5.37031796e+02, 9.79026534e-17
5.55904257e+02, 9.95926597e-17
5.75439937e+02, 1.01209847e-16
5.95662144e+02, 1.02754916e-16
6.16595002e+02, 1.04207158e-16
6.38263486e+02, 1.05573637e-16
6.60693448e+02, 1.06856509e-16
6.83911647e+02, 1.08055731e-16
7.07945784e+02, 1.09149640e-16
7.32824533e+02, 1.10139778e-16
7.58577575e+02, 1.11054500e-16
7.85235635e+02, 1.11861060e-16
8.12830516e+02, 1.12585065e-16
8.41395142e+02, 1.13205039e-16
8.70963590e+02, 1.13728628e-16
9.01571138e+02, 1.14155564e-16
9.33254301e+02, 1.14482614e-16
9.66050879e+02, 1.14734751e-16
1.00000000e+03, 1.14882647e-16
