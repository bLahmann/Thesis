1.00000000e+00, 9.88506890e-23
1.03514217e+00, 1.19861147e-22
1.07151931e+00, 1.45167858e-22
1.10917482e+00, 1.75299110e-22
1.14815362e+00, 2.11247150e-22
1.18850223e+00, 2.54285675e-22
1.23026877e+00, 3.04598756e-22
1.27350308e+00, 3.63777968e-22
1.31825674e+00, 4.34764267e-22
1.36458314e+00, 5.17474257e-22
1.41253754e+00, 6.14770092e-22
1.46217717e+00, 7.29878572e-22
1.51356125e+00, 8.63042132e-22
1.56675107e+00, 1.01726154e-21
1.62181010e+00, 1.19988822e-21
1.67880402e+00, 1.41219662e-21
1.73780083e+00, 1.65555222e-21
1.79887092e+00, 1.94128181e-21
1.86208714e+00, 2.26453842e-21
1.92752491e+00, 2.64370037e-21
1.99526231e+00, 3.07397209e-21
2.06538016e+00, 3.57321687e-21
2.13796209e+00, 4.14259679e-21
2.21309471e+00, 4.79316675e-21
2.29086765e+00, 5.53986590e-21
2.37137371e+00, 6.37589425e-21
2.45470892e+00, 7.34544443e-21
2.54097271e+00, 8.44584426e-21
2.63026799e+00, 9.67800706e-21
2.72270131e+00, 1.10843466e-20
2.81838293e+00, 1.26556699e-20
2.91742701e+00, 1.44535023e-20
3.01995172e+00, 1.64535725e-20
3.12607937e+00, 1.86947184e-20
3.23593657e+00, 2.12209624e-20
3.34965439e+00, 2.40489550e-20
3.46736850e+00, 2.72144462e-20
3.58921935e+00, 3.07325640e-20
3.71535229e+00, 3.46598356e-20
3.84591782e+00, 3.90410465e-20
3.98107171e+00, 4.38636207e-20
4.12097519e+00, 4.92616556e-20
4.26579519e+00, 5.52273874e-20
4.41570447e+00, 6.18266644e-20
4.57088190e+00, 6.90793702e-20
4.73151259e+00, 7.70859045e-20
4.89778819e+00, 8.59266676e-20
5.06990708e+00, 9.55644022e-20
5.24807460e+00, 1.06260500e-19
5.43250331e+00, 1.17989721e-19
5.62341325e+00, 1.30738919e-19
5.82103218e+00, 1.44766416e-19
6.02559586e+00, 1.60012730e-19
6.23734835e+00, 1.76721849e-19
6.45654229e+00, 1.94893267e-19
6.68343918e+00, 2.14541546e-19
6.91830971e+00, 2.36071376e-19
7.16143410e+00, 2.59371667e-19
7.41310241e+00, 2.84534970e-19
7.67361489e+00, 3.11952412e-19
7.94328235e+00, 3.41472916e-19
8.22242650e+00, 3.73186928e-19
8.51138038e+00, 4.07964083e-19
8.81048873e+00, 4.45127213e-19
9.12010839e+00, 4.84886606e-19
9.44060876e+00, 5.27841103e-19
9.77237221e+00, 5.74287316e-19
1.01157945e+01, 6.23830029e-19
1.04712855e+01, 6.77178649e-19
1.08392691e+01, 7.33846359e-19
1.12201845e+01, 7.95038661e-19
1.16144861e+01, 8.60088026e-19
1.20226443e+01, 9.29711001e-19
1.24451461e+01, 1.00389444e-18
1.28824955e+01, 1.08323010e-18
1.33352143e+01, 1.16736796e-18
1.38038426e+01, 1.25732737e-18
1.42889396e+01, 1.35237966e-18
1.47910839e+01, 1.45449641e-18
1.53108746e+01, 1.56200218e-18
1.58489319e+01, 1.67613161e-18
1.64058977e+01, 1.79656837e-18
1.69824365e+01, 1.92486383e-18
1.75792361e+01, 2.06015947e-18
1.81970086e+01, 2.20282995e-18
1.88364909e+01, 2.35480899e-18
1.94984460e+01, 2.51367392e-18
2.01836636e+01, 2.68245442e-18
2.08929613e+01, 2.86041753e-18
2.16271852e+01, 3.04663016e-18
2.23872114e+01, 3.24363672e-18
2.31739465e+01, 3.45048680e-18
2.39883292e+01, 3.66758442e-18
2.48313311e+01, 3.89711662e-18
2.57039578e+01, 4.13530041e-18
2.66072506e+01, 4.38871162e-18
2.75422870e+01, 4.65104972e-18
2.85101827e+01, 4.92808531e-18
2.95120923e+01, 5.21514031e-18
3.05492111e+01, 5.51798287e-18
3.16227766e+01, 5.83410933e-18
3.27340695e+01, 6.16409170e-18
3.38844156e+01, 6.50992022e-18
3.50751874e+01, 6.86967362e-18
3.63078055e+01, 7.24649276e-18
3.75837404e+01, 7.63748494e-18
3.89045145e+01, 8.04616318e-18
4.02717034e+01, 8.47294964e-18
4.16869383e+01, 8.91442386e-18
4.31519077e+01, 9.37389865e-18
4.46683592e+01, 9.85191142e-18
4.62381021e+01, 1.03492543e-17
4.78630092e+01, 1.08671124e-17
4.95450191e+01, 1.14014416e-17
5.12861384e+01, 1.19568087e-17
5.30884444e+01, 1.25338413e-17
5.49540874e+01, 1.31305870e-17
5.68852931e+01, 1.37485041e-17
5.88843655e+01, 1.43859029e-17
6.09536897e+01, 1.50479992e-17
6.30957344e+01, 1.57339158e-17
6.53130553e+01, 1.64399444e-17
6.76082975e+01, 1.71716875e-17
6.99841996e+01, 1.79263863e-17
7.24435960e+01, 1.87034356e-17
7.49894209e+01, 1.95052619e-17
7.76247117e+01, 2.03311546e-17
8.03526122e+01, 2.11821050e-17
8.31763771e+01, 2.20569773e-17
8.60993752e+01, 2.29614619e-17
8.91250938e+01, 2.38848323e-17
9.22571427e+01, 2.48407735e-17
9.54992586e+01, 2.58157851e-17
9.88553095e+01, 2.68292433e-17
1.02329299e+02, 2.78582012e-17
1.05925373e+02, 2.89193903e-17
1.09647820e+02, 3.00017781e-17
1.13501082e+02, 3.11139327e-17
1.17489755e+02, 3.22523125e-17
1.21618600e+02, 3.34186306e-17
1.25892541e+02, 3.46176534e-17
1.30316678e+02, 3.58331757e-17
1.34896288e+02, 3.70863032e-17
1.39636836e+02, 3.83651420e-17
1.44543977e+02, 3.96699526e-17
1.49623566e+02, 4.09992272e-17
1.54881662e+02, 4.23647055e-17
1.60324539e+02, 4.37563374e-17
1.65958691e+02, 4.51724702e-17
1.71790839e+02, 4.66240002e-17
1.77827941e+02, 4.81042595e-17
1.84077200e+02, 4.95919913e-17
1.90546072e+02, 5.11330557e-17
1.97242274e+02, 5.26935974e-17
2.04173794e+02, 5.42702823e-17
2.11348904e+02, 5.58869964e-17
2.18776162e+02, 5.75249368e-17
2.26464431e+02, 5.91986154e-17
2.34422882e+02, 6.08887418e-17
2.42661010e+02, 6.26101444e-17
2.51188643e+02, 6.43587756e-17
2.60015956e+02, 6.61390798e-17
2.69153480e+02, 6.79426681e-17
2.78612117e+02, 6.97706440e-17
2.88403150e+02, 7.16278188e-17
2.98538262e+02, 7.35039025e-17
3.09029543e+02, 7.53984053e-17
3.19889511e+02, 7.73357903e-17
3.31131121e+02, 7.92775418e-17
3.42767787e+02, 8.12608445e-17
3.54813389e+02, 8.32463165e-17
3.67282300e+02, 8.52603722e-17
3.80189396e+02, 8.73003506e-17
3.93550075e+02, 8.93532002e-17
4.07380278e+02, 9.14346993e-17
4.21696503e+02, 9.35330897e-17
4.36515832e+02, 9.56523266e-17
4.51855944e+02, 9.77748560e-17
4.67735141e+02, 9.99181907e-17
4.84172368e+02, 1.02070665e-16
5.01187234e+02, 1.04242652e-16
5.18800039e+02, 1.06437498e-16
5.37031796e+02, 1.08611636e-16
5.55904257e+02, 1.10811445e-16
5.75439937e+02, 1.13010350e-16
5.95662144e+02, 1.15197039e-16
6.16595002e+02, 1.17391477e-16
6.38263486e+02, 1.19585464e-16
6.60693448e+02, 1.21756207e-16
6.83911647e+02, 1.23912295e-16
7.07945784e+02, 1.26058260e-16
7.32824533e+02, 1.28175540e-16
7.58577575e+02, 1.30260120e-16
7.85235635e+02, 1.32298855e-16
8.12830516e+02, 1.34302980e-16
8.41395142e+02, 1.36256453e-16
8.70963590e+02, 1.38145355e-16
9.01571138e+02, 1.39978359e-16
9.33254301e+02, 1.41723443e-16
9.66050879e+02, 1.43397865e-16
1.00000000e+03, 1.44988322e-16
