1.00000000e+00, 2.69989898e-28
1.03514217e+00, 4.00136092e-28
1.07151931e+00, 5.70141257e-28
1.10917482e+00, 8.18058792e-28
1.14815362e+00, 1.14281704e-27
1.18850223e+00, 1.61793741e-27
1.23026877e+00, 2.34529700e-27
1.27350308e+00, 3.21245594e-27
1.31825674e+00, 4.48144453e-27
1.36458314e+00, 6.28624390e-27
1.41253754e+00, 8.77107136e-27
1.46217717e+00, 1.21613471e-26
1.51356125e+00, 1.68302031e-26
1.56675107e+00, 2.29631938e-26
1.62181010e+00, 3.20624482e-26
1.67880402e+00, 4.29722472e-26
1.73780083e+00, 5.80962048e-26
1.79887092e+00, 7.98238249e-26
1.86208714e+00, 1.05251667e-25
1.92752491e+00, 1.41551863e-25
1.99526231e+00, 1.89109082e-25
2.06538016e+00, 2.51107009e-25
2.13796209e+00, 3.34299009e-25
2.21309471e+00, 4.42295946e-25
2.29086765e+00, 5.84831807e-25
2.37137371e+00, 7.72225599e-25
2.45470892e+00, 1.00581466e-24
2.54097271e+00, 1.31377873e-24
2.63026799e+00, 1.72129544e-24
2.72270131e+00, 2.22098189e-24
2.81838293e+00, 2.84796510e-24
2.91742701e+00, 3.63268003e-24
3.01995172e+00, 4.72914823e-24
3.12607937e+00, 6.02611925e-24
3.23593657e+00, 7.69579886e-24
3.34965439e+00, 9.73279015e-24
3.46736850e+00, 1.24141461e-23
3.58921935e+00, 1.56841716e-23
3.71535229e+00, 1.96393366e-23
3.84591782e+00, 2.47733220e-23
3.98107171e+00, 3.11165957e-23
4.12097519e+00, 3.89263303e-23
4.26579519e+00, 4.82665138e-23
4.41570447e+00, 5.99853369e-23
4.57088190e+00, 7.44299603e-23
4.73151259e+00, 9.19813822e-23
4.89778819e+00, 1.12872848e-22
5.06990708e+00, 1.39286564e-22
5.24807460e+00, 1.69751993e-22
5.43250331e+00, 2.08065190e-22
5.62341325e+00, 2.52709913e-22
5.82103218e+00, 3.08114543e-22
6.02559586e+00, 3.74056478e-22
6.23734835e+00, 4.51602836e-22
6.45654229e+00, 5.43890570e-22
6.68343918e+00, 6.55583411e-22
6.91830971e+00, 7.86075739e-22
7.16143410e+00, 9.40613553e-22
7.41310241e+00, 1.12239896e-21
7.67361489e+00, 1.33940769e-21
7.94328235e+00, 1.59074189e-21
8.22242650e+00, 1.88651557e-21
8.51138038e+00, 2.23177522e-21
8.81048873e+00, 2.63105048e-21
9.12010839e+00, 3.10627048e-21
9.44060876e+00, 3.64323749e-21
9.77237221e+00, 4.27327444e-21
1.01157945e+01, 4.99681362e-21
1.04712855e+01, 5.82447351e-21
1.08392691e+01, 6.80081116e-21
1.12201845e+01, 7.88579571e-21
1.16144861e+01, 9.15617931e-21
1.20226443e+01, 1.05845036e-20
1.24451461e+01, 1.22392790e-20
1.28824955e+01, 1.41104938e-20
1.33352143e+01, 1.62177467e-20
1.38038426e+01, 1.86239268e-20
1.42889396e+01, 2.13369344e-20
1.47910839e+01, 2.43864994e-20
1.53108746e+01, 2.78156653e-20
1.58489319e+01, 3.17360477e-20
1.64058977e+01, 3.60146274e-20
1.69824365e+01, 4.08791918e-20
1.75792361e+01, 4.62590562e-20
1.81970086e+01, 5.23447588e-20
1.88364909e+01, 5.90703255e-20
1.94984460e+01, 6.65594681e-20
2.01836636e+01, 7.48324155e-20
2.08929613e+01, 8.39798993e-20
2.16271852e+01, 9.40382367e-20
2.23872114e+01, 1.05192020e-19
2.31739465e+01, 1.17456510e-19
2.39883292e+01, 1.30896847e-19
2.48313311e+01, 1.45703740e-19
2.57039578e+01, 1.61906569e-19
2.66072506e+01, 1.79491026e-19
2.75422870e+01, 1.98868234e-19
2.85101827e+01, 2.19931682e-19
2.95120923e+01, 2.42685824e-19
3.05492111e+01, 2.67405949e-19
3.16227766e+01, 2.94422820e-19
3.27340695e+01, 3.23349407e-19
3.38844156e+01, 3.54773642e-19
3.50751874e+01, 3.88969737e-19
3.63078055e+01, 4.25348562e-19
3.75837404e+01, 4.64668923e-19
3.89045145e+01, 5.06985354e-19
4.02717034e+01, 5.52380412e-19
4.16869383e+01, 6.00801979e-19
4.31519077e+01, 6.52872809e-19
4.46683592e+01, 7.08430463e-19
4.62381021e+01, 7.67824204e-19
4.78630092e+01, 8.30767321e-19
4.95450191e+01, 8.97744423e-19
5.12861384e+01, 9.69101800e-19
5.30884444e+01, 1.04516201e-18
5.49540874e+01, 1.12577368e-18
5.68852931e+01, 1.21008774e-18
5.88843655e+01, 1.30017726e-18
6.09536897e+01, 1.39522961e-18
6.30957344e+01, 1.49535643e-18
6.53130553e+01, 1.60083769e-18
6.76082975e+01, 1.71198049e-18
6.99841996e+01, 1.82959577e-18
7.24435960e+01, 1.95150182e-18
7.49894209e+01, 2.08034773e-18
7.76247117e+01, 2.21521593e-18
8.03526122e+01, 2.35568005e-18
8.31763771e+01, 2.50422142e-18
8.60993752e+01, 2.65774955e-18
8.91250938e+01, 2.81935161e-18
9.22571427e+01, 2.98626481e-18
9.54992586e+01, 3.16123789e-18
9.88553095e+01, 3.34190586e-18
1.02329299e+02, 3.52986640e-18
1.05925373e+02, 3.72650272e-18
1.09647820e+02, 3.92943698e-18
1.13501082e+02, 4.13964573e-18
1.17489755e+02, 4.35682892e-18
1.21618600e+02, 4.58221793e-18
1.25892541e+02, 4.81313875e-18
1.30316678e+02, 5.05370417e-18
1.34896288e+02, 5.29930699e-18
1.39636836e+02, 5.55254760e-18
1.44543977e+02, 5.81554740e-18
1.49623566e+02, 6.08267544e-18
1.54881662e+02, 6.35826895e-18
1.60324539e+02, 6.64228121e-18
1.65958691e+02, 6.93040365e-18
1.71790839e+02, 7.22504899e-18
1.77827941e+02, 7.53014601e-18
1.84077200e+02, 7.84049517e-18
1.90546072e+02, 8.15453355e-18
1.97242274e+02, 8.47571422e-18
2.04173794e+02, 8.80253731e-18
2.11348904e+02, 9.13649287e-18
2.18776162e+02, 9.47657667e-18
2.26464431e+02, 9.82070619e-18
2.34422882e+02, 1.01695914e-17
2.42661010e+02, 1.05240320e-17
2.51188643e+02, 1.08837075e-17
2.60015956e+02, 1.12460802e-17
2.69153480e+02, 1.16156776e-17
2.78612117e+02, 1.19861108e-17
2.88403150e+02, 1.23627630e-17
2.98538262e+02, 1.27428742e-17
3.09029543e+02, 1.31253109e-17
3.19889511e+02, 1.35119102e-17
3.31131121e+02, 1.39048301e-17
3.42767787e+02, 1.42971833e-17
3.54813389e+02, 1.46951745e-17
3.67282300e+02, 1.50952395e-17
3.80189396e+02, 1.55001316e-17
3.93550075e+02, 1.59092492e-17
4.07380278e+02, 1.63168935e-17
4.21696503e+02, 1.67346459e-17
4.36515832e+02, 1.71532684e-17
4.51855944e+02, 1.75755020e-17
4.67735141e+02, 1.80031571e-17
4.84172368e+02, 1.84355139e-17
5.01187234e+02, 1.88728332e-17
5.18800039e+02, 1.93145980e-17
5.37031796e+02, 1.97618159e-17
5.55904257e+02, 2.02153377e-17
5.75439937e+02, 2.06796269e-17
5.95662144e+02, 2.11473409e-17
6.16595002e+02, 2.16265865e-17
6.38263486e+02, 2.21125320e-17
6.60693448e+02, 2.26071293e-17
6.83911647e+02, 2.31093311e-17
7.07945784e+02, 2.36270452e-17
7.32824533e+02, 2.41523396e-17
7.58577575e+02, 2.46933525e-17
7.85235635e+02, 2.52416575e-17
8.12830516e+02, 2.58076263e-17
8.41395142e+02, 2.63845082e-17
8.70963590e+02, 2.69813651e-17
9.01571138e+02, 2.75918394e-17
9.33254301e+02, 2.82185426e-17
9.66050879e+02, 2.88550633e-17
1.00000000e+03, 2.95191168e-17
