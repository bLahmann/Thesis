1.00000000e+00, 3.62065259e-26
1.03514217e+00, 5.02425922e-26
1.07151931e+00, 7.20329992e-26
1.10917482e+00, 9.93162190e-26
1.14815362e+00, 1.35987694e-25
1.18850223e+00, 1.91908640e-25
1.23026877e+00, 2.63280179e-25
1.27350308e+00, 3.61714224e-25
1.31825674e+00, 4.92071128e-25
1.36458314e+00, 6.80240004e-25
1.41253754e+00, 9.09933756e-25
1.46217717e+00, 1.23187708e-24
1.51356125e+00, 1.69267040e-24
1.56675107e+00, 2.24820241e-24
1.62181010e+00, 2.99845660e-24
1.67880402e+00, 3.98756292e-24
1.73780083e+00, 5.30803427e-24
1.79887092e+00, 7.06824946e-24
1.86208714e+00, 9.30286589e-24
1.92752491e+00, 1.21036167e-23
1.99526231e+00, 1.60075712e-23
2.06538016e+00, 2.10302542e-23
2.13796209e+00, 2.73848601e-23
2.21309471e+00, 3.54332229e-23
2.29086765e+00, 4.56477063e-23
2.37137371e+00, 5.91438407e-23
2.45470892e+00, 7.56767531e-23
2.54097271e+00, 9.71782145e-23
2.63026799e+00, 1.24676890e-22
2.72270131e+00, 1.58694458e-22
2.81838293e+00, 2.01459414e-22
2.91742701e+00, 2.55807074e-22
3.01995172e+00, 3.24352531e-22
3.12607937e+00, 4.07659983e-22
3.23593657e+00, 5.15039919e-22
3.34965439e+00, 6.41171400e-22
3.46736850e+00, 8.04089239e-22
3.58921935e+00, 9.96710902e-22
3.71535229e+00, 1.24710088e-21
3.84591782e+00, 1.54578134e-21
3.98107171e+00, 1.90213735e-21
4.12097519e+00, 2.35370523e-21
4.26579519e+00, 2.89429245e-21
4.41570447e+00, 3.55259857e-21
4.57088190e+00, 4.35035279e-21
4.73151259e+00, 5.30812525e-21
4.89778819e+00, 6.49623364e-21
5.06990708e+00, 7.88544516e-21
5.24807460e+00, 9.56587510e-21
5.43250331e+00, 1.15949468e-20
5.62341325e+00, 1.39708500e-20
5.82103218e+00, 1.68523434e-20
6.02559586e+00, 2.02925443e-20
6.23734835e+00, 2.43085278e-20
6.45654229e+00, 2.91006820e-20
6.68343918e+00, 3.47744927e-20
6.91830971e+00, 4.15555759e-20
7.16143410e+00, 4.93783240e-20
7.41310241e+00, 5.85992501e-20
7.67361489e+00, 6.96463034e-20
7.94328235e+00, 8.23951183e-20
8.22242650e+00, 9.72673057e-20
8.51138038e+00, 1.14586663e-19
8.81048873e+00, 1.35071144e-19
9.12010839e+00, 1.58460943e-19
9.44060876e+00, 1.85801834e-19
9.77237221e+00, 2.17872205e-19
1.01157945e+01, 2.54484516e-19
1.04712855e+01, 2.96967925e-19
1.08392691e+01, 3.46507576e-19
1.12201845e+01, 4.02712936e-19
1.16144861e+01, 4.67506078e-19
1.20226443e+01, 5.42069190e-19
1.24451461e+01, 6.28089020e-19
1.28824955e+01, 7.26349671e-19
1.33352143e+01, 8.38228781e-19
1.38038426e+01, 9.66929539e-19
1.42889396e+01, 1.11216972e-18
1.47910839e+01, 1.27963208e-18
1.53108746e+01, 1.46775585e-18
1.58489319e+01, 1.68415337e-18
1.64058977e+01, 1.92655543e-18
1.69824365e+01, 2.20298044e-18
1.75792361e+01, 2.51224183e-18
1.81970086e+01, 2.86449081e-18
1.88364909e+01, 3.25780991e-18
1.94984460e+01, 3.70276316e-18
2.01836636e+01, 4.20556181e-18
2.08929613e+01, 4.76032755e-18
2.16271852e+01, 5.38403609e-18
2.23872114e+01, 6.07887707e-18
2.31739465e+01, 6.85571861e-18
2.39883292e+01, 7.71461930e-18
2.48313311e+01, 8.67578078e-18
2.57039578e+01, 9.72688587e-18
2.66072506e+01, 1.08826748e-17
2.75422870e+01, 1.21702328e-17
2.85101827e+01, 1.35793060e-17
2.95120923e+01, 1.51203586e-17
3.05492111e+01, 1.68052396e-17
3.16227766e+01, 1.86420681e-17
3.27340695e+01, 2.06279690e-17
3.38844156e+01, 2.27830411e-17
3.50751874e+01, 2.51494294e-17
3.63078055e+01, 2.76476353e-17
3.75837404e+01, 3.03616491e-17
3.89045145e+01, 3.32663740e-17
4.02717034e+01, 3.63752112e-17
4.16869383e+01, 3.96869236e-17
4.31519077e+01, 4.31849306e-17
4.46683592e+01, 4.69199320e-17
4.62381021e+01, 5.08622635e-17
4.78630092e+01, 5.49901130e-17
4.95450191e+01, 5.93280579e-17
5.12861384e+01, 6.39121985e-17
5.30884444e+01, 6.86977695e-17
5.49540874e+01, 7.36317892e-17
5.68852931e+01, 7.87634938e-17
5.88843655e+01, 8.40872051e-17
6.09536897e+01, 8.96310571e-17
6.30957344e+01, 9.52397879e-17
6.53130553e+01, 1.01056551e-16
6.76082975e+01, 1.06988596e-16
6.99841996e+01, 1.13072356e-16
7.24435960e+01, 1.19196491e-16
7.49894209e+01, 1.25465467e-16
7.76247117e+01, 1.31714151e-16
8.03526122e+01, 1.38082459e-16
8.31763771e+01, 1.44446404e-16
8.60993752e+01, 1.50845418e-16
8.91250938e+01, 1.57190841e-16
9.22571427e+01, 1.63590184e-16
9.54992586e+01, 1.69857170e-16
9.88553095e+01, 1.76074685e-16
1.02329299e+02, 1.82220401e-16
1.05925373e+02, 1.88216064e-16
1.09647820e+02, 1.94114670e-16
1.13501082e+02, 1.99843263e-16
1.17489755e+02, 2.05410500e-16
1.21618600e+02, 2.10783012e-16
1.25892541e+02, 2.15986532e-16
1.30316678e+02, 2.20958562e-16
1.34896288e+02, 2.25653438e-16
1.39636836e+02, 2.30141410e-16
1.44543977e+02, 2.34367147e-16
1.49623566e+02, 2.38256267e-16
1.54881662e+02, 2.41900813e-16
1.60324539e+02, 2.45281965e-16
1.65958691e+02, 2.48298880e-16
1.71790839e+02, 2.51020828e-16
1.77827941e+02, 2.53445127e-16
1.84077200e+02, 2.55530644e-16
1.90546072e+02, 2.57271819e-16
1.97242274e+02, 2.58702037e-16
2.04173794e+02, 2.59789338e-16
2.11348904e+02, 2.60517506e-16
2.18776162e+02, 2.60976693e-16
2.26464431e+02, 2.61112832e-16
2.34422882e+02, 2.60878993e-16
2.42661010e+02, 2.60352594e-16
2.51188643e+02, 2.59476573e-16
2.60015956e+02, 2.58357274e-16
2.69153480e+02, 2.56907672e-16
2.78612117e+02, 2.55151363e-16
2.88403150e+02, 2.53128437e-16
2.98538262e+02, 2.50853143e-16
3.09029543e+02, 2.48341864e-16
3.19889511e+02, 2.45616353e-16
3.31131121e+02, 2.42595461e-16
3.42767787e+02, 2.39396672e-16
3.54813389e+02, 2.35994606e-16
3.67282300e+02, 2.32383328e-16
3.80189396e+02, 2.28708048e-16
3.93550075e+02, 2.24753869e-16
4.07380278e+02, 2.20742428e-16
4.21696503e+02, 2.16515530e-16
4.36515832e+02, 2.12271720e-16
4.51855944e+02, 2.07858674e-16
4.67735141e+02, 2.03424972e-16
4.84172368e+02, 1.98841642e-16
5.01187234e+02, 1.94217250e-16
5.18800039e+02, 1.89597293e-16
5.37031796e+02, 1.84907327e-16
5.55904257e+02, 1.80137339e-16
5.75439937e+02, 1.75472312e-16
5.95662144e+02, 1.70695601e-16
6.16595002e+02, 1.66001872e-16
6.38263486e+02, 1.61267505e-16
6.60693448e+02, 1.56611560e-16
6.83911647e+02, 1.51946493e-16
7.07945784e+02, 1.47345105e-16
7.32824533e+02, 1.42811849e-16
7.58577575e+02, 1.38302234e-16
7.85235635e+02, 1.33871532e-16
8.12830516e+02, 1.29492990e-16
8.41395142e+02, 1.25167944e-16
8.70963590e+02, 1.20983210e-16
9.01571138e+02, 1.16803570e-16
9.33254301e+02, 1.12770723e-16
9.66050879e+02, 1.08794441e-16
1.00000000e+03, 1.04881428e-16
