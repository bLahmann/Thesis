1.00000000e+00, 3.97061096e-37
1.03514217e+00, 1.74178792e-30
1.07151931e+00, 2.87950990e-31
1.10917482e+00, 2.57932674e-31
1.14815362e+00, 4.79615662e-30
1.18850223e+00, 1.30673795e-31
1.23026877e+00, 4.97357705e-30
1.27350308e+00, 1.01526356e-29
1.31825674e+00, 1.87673465e-29
1.36458314e+00, 3.40255726e-29
1.41253754e+00, 5.30775050e-29
1.46217717e+00, 6.97593915e-29
1.51356125e+00, 1.63051398e-28
1.56675107e+00, 2.25834688e-28
1.62181010e+00, 3.02153720e-28
1.67880402e+00, 4.89223738e-28
1.73780083e+00, 7.43298210e-28
1.79887092e+00, 1.05779410e-27
1.86208714e+00, 1.42284958e-27
1.92752491e+00, 2.03123652e-27
1.99526231e+00, 2.88466167e-27
2.06538016e+00, 4.06611056e-27
2.13796209e+00, 5.67033059e-27
2.21309471e+00, 7.82403072e-27
2.29086765e+00, 1.09669995e-26
2.37137371e+00, 1.40280582e-26
2.45470892e+00, 1.90304366e-26
2.54097271e+00, 2.52561109e-26
2.63026799e+00, 3.27101900e-26
2.72270131e+00, 4.32124038e-26
2.81838293e+00, 5.56684574e-26
2.91742701e+00, 7.13073569e-26
3.01995172e+00, 9.04175279e-26
3.12607937e+00, 1.19278500e-25
3.23593657e+00, 1.46421554e-25
3.34965439e+00, 1.89162135e-25
3.46736850e+00, 2.46525296e-25
3.58921935e+00, 3.39749080e-25
3.71535229e+00, 4.10133119e-25
3.84591782e+00, 5.12175856e-25
3.98107171e+00, 6.58751205e-25
4.12097519e+00, 8.84118991e-25
4.26579519e+00, 1.17028916e-24
4.41570447e+00, 1.45811530e-24
4.57088190e+00, 1.85873421e-24
4.73151259e+00, 2.45956600e-24
4.89778819e+00, 3.24798758e-24
5.06990708e+00, 4.27004278e-24
5.24807460e+00, 5.60462138e-24
5.43250331e+00, 7.43825064e-24
5.62341325e+00, 9.52759859e-24
5.82103218e+00, 1.25042547e-23
6.02559586e+00, 1.66998144e-23
6.23734835e+00, 2.10114059e-23
6.45654229e+00, 2.78997605e-23
6.68343918e+00, 3.62516973e-23
6.91830971e+00, 4.71215414e-23
7.16143410e+00, 5.80149210e-23
7.41310241e+00, 7.42611312e-23
7.67361489e+00, 9.30667414e-23
7.94328235e+00, 1.21942988e-22
8.22242650e+00, 1.54436825e-22
8.51138038e+00, 1.92064077e-22
8.81048873e+00, 2.48991806e-22
9.12010839e+00, 3.07431846e-22
9.44060876e+00, 3.98433666e-22
9.77237221e+00, 4.91809669e-22
1.01157945e+01, 6.06791776e-22
1.04712855e+01, 7.58921229e-22
1.08392691e+01, 9.61896471e-22
1.12201845e+01, 1.21309063e-21
1.16144861e+01, 1.49730484e-21
1.20226443e+01, 1.87435977e-21
1.24451461e+01, 2.32797650e-21
1.28824955e+01, 2.88851065e-21
1.33352143e+01, 3.52448549e-21
1.38038426e+01, 4.40744745e-21
1.42889396e+01, 5.44485666e-21
1.47910839e+01, 6.78958205e-21
1.53108746e+01, 8.21379540e-21
1.58489319e+01, 1.00554878e-20
1.64058977e+01, 1.21468158e-20
1.69824365e+01, 1.48010526e-20
1.75792361e+01, 1.80615601e-20
1.81970086e+01, 2.17544693e-20
1.88364909e+01, 2.63548082e-20
1.94984460e+01, 3.15459674e-20
2.01836636e+01, 3.81185859e-20
2.08929613e+01, 4.55489100e-20
2.16271852e+01, 5.40757151e-20
2.23872114e+01, 6.46782797e-20
2.31739465e+01, 7.71202621e-20
2.39883292e+01, 9.17299658e-20
2.48313311e+01, 1.08711773e-19
2.57039578e+01, 1.28472467e-19
2.66072506e+01, 1.51818581e-19
2.75422870e+01, 1.80551156e-19
2.85101827e+01, 2.11262732e-19
2.95120923e+01, 2.47928722e-19
3.05492111e+01, 2.90415817e-19
3.16227766e+01, 3.43333428e-19
3.27340695e+01, 3.99583108e-19
3.38844156e+01, 4.70446541e-19
3.50751874e+01, 5.44593875e-19
3.63078055e+01, 6.32207146e-19
3.75837404e+01, 7.33724859e-19
3.89045145e+01, 8.48971298e-19
4.02717034e+01, 9.82872175e-19
4.16869383e+01, 1.13399502e-18
4.31519077e+01, 1.30188175e-18
4.46683592e+01, 1.49412759e-18
4.62381021e+01, 1.71911666e-18
4.78630092e+01, 1.96271613e-18
4.95450191e+01, 2.22985867e-18
5.12861384e+01, 2.52921103e-18
5.30884444e+01, 2.88095342e-18
5.49540874e+01, 3.26424754e-18
5.68852931e+01, 3.68977585e-18
5.88843655e+01, 4.15230206e-18
6.09536897e+01, 4.66813545e-18
6.30957344e+01, 5.25024167e-18
6.53130553e+01, 5.86887344e-18
6.76082975e+01, 6.56115912e-18
6.99841996e+01, 7.31837011e-18
7.24435960e+01, 8.15060535e-18
7.49894209e+01, 9.03976290e-18
7.76247117e+01, 1.00542979e-17
8.03526122e+01, 1.11096724e-17
8.31763771e+01, 1.22279519e-17
8.60993752e+01, 1.34927679e-17
8.91250938e+01, 1.48897688e-17
9.22571427e+01, 1.63190050e-17
9.54992586e+01, 1.78684047e-17
9.88553095e+01, 1.95603479e-17
1.02329299e+02, 2.13347030e-17
1.05925373e+02, 2.32797743e-17
1.09647820e+02, 2.53287650e-17
1.13501082e+02, 2.75532986e-17
1.17489755e+02, 2.98739948e-17
1.21618600e+02, 3.23667607e-17
1.25892541e+02, 3.50283798e-17
1.30316678e+02, 3.78196235e-17
1.34896288e+02, 4.07670303e-17
1.39636836e+02, 4.39150802e-17
1.44543977e+02, 4.72330757e-17
1.49623566e+02, 5.07741784e-17
1.54881662e+02, 5.44513527e-17
1.60324539e+02, 5.82961193e-17
1.65958691e+02, 6.24129909e-17
1.71790839e+02, 6.65775343e-17
1.77827941e+02, 7.11078488e-17
1.84077200e+02, 7.56857813e-17
1.90546072e+02, 8.05122843e-17
1.97242274e+02, 8.57534745e-17
2.04173794e+02, 9.09001106e-17
2.11348904e+02, 9.63518899e-17
2.18776162e+02, 1.02026402e-16
2.26464431e+02, 1.07929511e-16
2.34422882e+02, 1.14048334e-16
2.42661010e+02, 1.20345279e-16
2.51188643e+02, 1.26834427e-16
2.60015956e+02, 1.33643547e-16
2.69153480e+02, 1.40389083e-16
2.78612117e+02, 1.47590767e-16
2.88403150e+02, 1.54973572e-16
2.98538262e+02, 1.62311869e-16
3.09029543e+02, 1.69990114e-16
3.19889511e+02, 1.77878058e-16
3.31131121e+02, 1.86147573e-16
3.42767787e+02, 1.94282784e-16
3.54813389e+02, 2.02611692e-16
3.67282300e+02, 2.11299027e-16
3.80189396e+02, 2.20265399e-16
3.93550075e+02, 2.29301119e-16
4.07380278e+02, 2.38307575e-16
4.21696503e+02, 2.47622476e-16
4.36515832e+02, 2.56897531e-16
4.51855944e+02, 2.66791543e-16
4.67735141e+02, 2.76523743e-16
4.84172368e+02, 2.86497116e-16
5.01187234e+02, 2.96538154e-16
5.18800039e+02, 3.06663023e-16
5.37031796e+02, 3.16941715e-16
5.55904257e+02, 3.27509616e-16
5.75439937e+02, 3.37932447e-16
5.95662144e+02, 3.48790355e-16
6.16595002e+02, 3.59366267e-16
6.38263486e+02, 3.70750627e-16
6.60693448e+02, 3.81435735e-16
6.83911647e+02, 3.92651300e-16
7.07945784e+02, 4.03605670e-16
7.32824533e+02, 4.15431344e-16
7.58577575e+02, 4.27051427e-16
7.85235635e+02, 4.38437326e-16
8.12830516e+02, 4.49944934e-16
8.41395142e+02, 4.61715256e-16
8.70963590e+02, 4.73405763e-16
9.01571138e+02, 4.85026676e-16
9.33254301e+02, 4.97021958e-16
9.66050879e+02, 5.09192129e-16
1.00000000e+03, 5.21196355e-16
